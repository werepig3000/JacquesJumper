library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity crouchFinalROM is

  port(

  clk : in std_logic;
  x_address: in unsigned(4 downto 0); 
  y_address: in unsigned(5 downto 0);
  rgb : out std_logic_vector(5 downto 0)

      );

end crouchFinalROM;


architecture synth of crouchFinalROM is

signal xy_address : std_logic_vector(10 downto 0); 


begin

   process (clk) begin

if rising_edge(clk) then

case xy_address is


when "01110101011" => rgb <= "101010";
when "01110110001" => rgb <= "101010";
when "01110110010" => rgb <= "101010";
when "01111001001" => rgb <= "100101";
when "01111001010" => rgb <= "111001";
when "01111001011" => rgb <= "011001";
when "01111001100" => rgb <= "101010";
when "01111001101" => rgb <= "101010";
when "01111001110" => rgb <= "101010";
when "01111001111" => rgb <= "101010";
when "01111010000" => rgb <= "101010";
when "01111010001" => rgb <= "010101";
when "01111010010" => rgb <= "111001";
when "01111010011" => rgb <= "010101";
when "01111101001" => rgb <= "010000";
when "01111101010" => rgb <= "111000";
when "01111101011" => rgb <= "010100";
when "01111101100" => rgb <= "011001";
when "01111101101" => rgb <= "011001";
when "01111101110" => rgb <= "101001";
when "01111101111" => rgb <= "011001";
when "01111110000" => rgb <= "011000";
when "01111110001" => rgb <= "010100";
when "01111110010" => rgb <= "101000";
when "01111110011" => rgb <= "111001";
when "10000001001" => rgb <= "101001";
when "10000001010" => rgb <= "101000";
when "10000001011" => rgb <= "011001";
when "10000001100" => rgb <= "011001";
when "10000001101" => rgb <= "100100";
when "10000001110" => rgb <= "100100";
when "10000001111" => rgb <= "100100";
when "10000010000" => rgb <= "011000";
when "10000010001" => rgb <= "011001";
when "10000010010" => rgb <= "100100";
when "10000010011" => rgb <= "111001";
when "10000101010" => rgb <= "101010";
when "10000101011" => rgb <= "101001";
when "10000101100" => rgb <= "100101";
when "10000101101" => rgb <= "100101";
when "10000101110" => rgb <= "100101";
when "10000101111" => rgb <= "100101";
when "10000110000" => rgb <= "100101";
when "10000110001" => rgb <= "100101";
when "10000110010" => rgb <= "011001";
when "10000110011" => rgb <= "101001";
when "10001001011" => rgb <= "101010";
when "10001001100" => rgb <= "101010";
when "10001001101" => rgb <= "101010";
when "10001001110" => rgb <= "101010";
when "10001001111" => rgb <= "101010";
when "10001010000" => rgb <= "101010";
when "10001010001" => rgb <= "101010";
when "10001010010" => rgb <= "101010";
when "10001101011" => rgb <= "101010";
when "10001101100" => rgb <= "101010";
when "10001101101" => rgb <= "101010";
when "10001101110" => rgb <= "101010";
when "10001101111" => rgb <= "101010";
when "10001110000" => rgb <= "101010";
when "10001110001" => rgb <= "101010";
when "10001110010" => rgb <= "101010";
when "10010001010" => rgb <= "101010";
when "10010001011" => rgb <= "101010";
when "10010001100" => rgb <= "101010";
when "10010001101" => rgb <= "101010";
when "10010001110" => rgb <= "101010";
when "10010001111" => rgb <= "101010";
when "10010010000" => rgb <= "101010";
when "10010010001" => rgb <= "101010";
when "10010010010" => rgb <= "101010";
when "10010101001" => rgb <= "010101";
when "10010101010" => rgb <= "101010";
when "10010101011" => rgb <= "101001";
when "10010101100" => rgb <= "101010";
when "10010101101" => rgb <= "101010";
when "10010101110" => rgb <= "101010";
when "10010101111" => rgb <= "101010";
when "10010110000" => rgb <= "101010";
when "10010110001" => rgb <= "101010";
when "10010110010" => rgb <= "101010";
when "10010110011" => rgb <= "100101";
when "10011001000" => rgb <= "010101";
when "10011001001" => rgb <= "101010";
when "10011001010" => rgb <= "100011";
when "10011001011" => rgb <= "100101";
when "10011001100" => rgb <= "101010";
when "10011001101" => rgb <= "101010";
when "10011001110" => rgb <= "101010";
when "10011001111" => rgb <= "101010";
when "10011010000" => rgb <= "101010";
when "10011010001" => rgb <= "101010";
when "10011010010" => rgb <= "100011";
when "10011010011" => rgb <= "101010";
when "10011010100" => rgb <= "010101";
when "10011010101" => rgb <= "010101";
when "10011010110" => rgb <= "101010";
when "10011100011" => rgb <= "010101";
when "10011100100" => rgb <= "010101";
when "10011100101" => rgb <= "010101";
when "10011100110" => rgb <= "010101";
when "10011100111" => rgb <= "010101";
when "10011101000" => rgb <= "100101";
when "10011101001" => rgb <= "010101";
when "10011101010" => rgb <= "010101";
when "10011101011" => rgb <= "010101";
when "10011101100" => rgb <= "101010";
when "10011101101" => rgb <= "101010";
when "10011101110" => rgb <= "101001";
when "10011101111" => rgb <= "101001";
when "10011110000" => rgb <= "101010";
when "10011110001" => rgb <= "100101";
when "10011110010" => rgb <= "101010";
when "10011110011" => rgb <= "101001";
when "10011110100" => rgb <= "010101";
when "10011110101" => rgb <= "010101";
when "10011110110" => rgb <= "010100";
when "10011110111" => rgb <= "010101";
when "10011111000" => rgb <= "010101";
when "10100000101" => rgb <= "010101";
when "10100000110" => rgb <= "010101";
when "10100000111" => rgb <= "010101";
when "10100001000" => rgb <= "010101";
when "10100001001" => rgb <= "010101";
when "10100001010" => rgb <= "010101";
when "10100001011" => rgb <= "010101";
when "10100001100" => rgb <= "010101";
when "10100001101" => rgb <= "101001";
when "10100001110" => rgb <= "101001";
when "10100001111" => rgb <= "101001";
when "10100010000" => rgb <= "100101";
when "10100010001" => rgb <= "010101";
when "10100010010" => rgb <= "010101";
when "10100010011" => rgb <= "010101";
when "10100010100" => rgb <= "010101";
when "10100010101" => rgb <= "100101";
when "10100010110" => rgb <= "011001";
when "10100010111" => rgb <= "010101";
when "10100011000" => rgb <= "010101";
when "10100100101" => rgb <= "100101";
when "10100100110" => rgb <= "100101";
when "10100100111" => rgb <= "100101";
when "10100101001" => rgb <= "100101";
when "10100101010" => rgb <= "100101";
when "10100101011" => rgb <= "010101";
when "10100101100" => rgb <= "010101";
when "10100101101" => rgb <= "010101";
when "10100101110" => rgb <= "100101";
when "10100101111" => rgb <= "010101";
when "10100110000" => rgb <= "010101";
when "10100110001" => rgb <= "010101";
when "10100110010" => rgb <= "010101";
when "10100110011" => rgb <= "010101";
when "10100110100" => rgb <= "010101";
when "10100110101" => rgb <= "100101";
when "10100110110" => rgb <= "010100";
when "10100110111" => rgb <= "010101";
when "10101000010" => rgb <= "101010";
when "10101000011" => rgb <= "100101";
when "10101000100" => rgb <= "100101";
when "10101000101" => rgb <= "100101";
when "10101000110" => rgb <= "100101";
when "10101000111" => rgb <= "101010";
when "10101001100" => rgb <= "010110";
when "10101001101" => rgb <= "010101";
when "10101001110" => rgb <= "010101";
when "10101001111" => rgb <= "010101";
when "10101010000" => rgb <= "010101";
when "10101010001" => rgb <= "010101";
when "10101010110" => rgb <= "010100";
when "10101010111" => rgb <= "010100";
when "10101011000" => rgb <= "010101";
when "10101011001" => rgb <= "100101";
when "10101100000" => rgb <= "100101";
when "10101100001" => rgb <= "100101";
when "10101100010" => rgb <= "100101";
when "10101100011" => rgb <= "100101";
when "10101100100" => rgb <= "100101";
when "10101100101" => rgb <= "100101";
when "10101100111" => rgb <= "101001";
when "10101110110" => rgb <= "010101";
when "10101110111" => rgb <= "100101";
when "10101111001" => rgb <= "100101";
when "10101111010" => rgb <= "100101";
when "10110000010" => rgb <= "100101";
when "10110000101" => rgb <= "101010";
when "10110000110" => rgb <= "100101";
when "10110000111" => rgb <= "100101";
when "10110001000" => rgb <= "100101";
when "10110001001" => rgb <= "100101";
when "10110001010" => rgb <= "100101";
when "10110010101" => rgb <= "100101";
when "10110010110" => rgb <= "100101";
when "10110010111" => rgb <= "101001";
when "10110100011" => rgb <= "100101";
when "10110100100" => rgb <= "101010";
when "10110100101" => rgb <= "101010";
when "10110100111" => rgb <= "101001";
when "10110110011" => rgb <= "100101";
when "10110110100" => rgb <= "100101";
when "10110110101" => rgb <= "100101";
when "10110110110" => rgb <= "100101";
when "10110111001" => rgb <= "101001";
when "10110111010" => rgb <= "100101";
when "10111000111" => rgb <= "101010";
when "10111010101" => rgb <= "100101";
when others => rgb <= "110011";




end case;

end if;

   end process;

   xy_address <= std_logic_vector(y_address) & std_logic_vector(x_address);
   
end;