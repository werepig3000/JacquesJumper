library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity crouch1ROM is

  port(

  clk : in std_logic;
  x_address: in unsigned(4 downto 0); 
  y_address: in unsigned(5 downto 0);
  rgb : out std_logic_vector(5 downto 0)

      );

end crouch1ROM;


architecture synth of crouch1ROM is

signal xy_address : std_logic_vector(10 downto 0); 


begin

   process (clk) begin

if rising_edge(clk) then

case xy_address is


when "00001101010" => rgb <= "101010";
when "00001101011" => rgb <= "101010";
when "00001101100" => rgb <= "101110";
when "00001101101" => rgb <= "101110";
when "00001101110" => rgb <= "101010";
when "00001101111" => rgb <= "101010";
when "00010001010" => rgb <= "010101";
when "00010001011" => rgb <= "011001";
when "00010001100" => rgb <= "101110";
when "00010001101" => rgb <= "101110";
when "00010001110" => rgb <= "011001";
when "00010001111" => rgb <= "100101";
when "00010101010" => rgb <= "010100";
when "00010101011" => rgb <= "011001";
when "00010101100" => rgb <= "101110";
when "00010101101" => rgb <= "101101";
when "00010101110" => rgb <= "011001";
when "00010101111" => rgb <= "010100";
when "00011001010" => rgb <= "010101";
when "00011001011" => rgb <= "011001";
when "00011001100" => rgb <= "011001";
when "00011001101" => rgb <= "101101";
when "00011001110" => rgb <= "011001";
when "00011001111" => rgb <= "010100";
when "00011101001" => rgb <= "101010";
when "00011101010" => rgb <= "011001";
when "00011101011" => rgb <= "011001";
when "00011101100" => rgb <= "011001";
when "00011101101" => rgb <= "011000";
when "00011101110" => rgb <= "010100";
when "00011101111" => rgb <= "010100";
when "00100001010" => rgb <= "101001";
when "00100001011" => rgb <= "011001";
when "00100001100" => rgb <= "011001";
when "00100001101" => rgb <= "010101";
when "00100001110" => rgb <= "010101";
when "00100001111" => rgb <= "010101";
when "00100101010" => rgb <= "101010";
when "00100101011" => rgb <= "101001";
when "00100101100" => rgb <= "011001";
when "00100101101" => rgb <= "010101";
when "00100101110" => rgb <= "010101";
when "00100101111" => rgb <= "010101";
when "00101001010" => rgb <= "101010";
when "00101001011" => rgb <= "101001";
when "00101001100" => rgb <= "011001";
when "00101001101" => rgb <= "010101";
when "00101001110" => rgb <= "010101";
when "00101001111" => rgb <= "010101";
when "00101101010" => rgb <= "011001";
when "00101101011" => rgb <= "101001";
when "00101101100" => rgb <= "011001";
when "00101101101" => rgb <= "010101";
when "00101101110" => rgb <= "010101";
when "00101101111" => rgb <= "010101";
when "00101110000" => rgb <= "010101";
when "00101110001" => rgb <= "101010";
when "00110001001" => rgb <= "011001";
when "00110001010" => rgb <= "010101";
when "00110001011" => rgb <= "010101";
when "00110001100" => rgb <= "101001";
when "00110001101" => rgb <= "010101";
when "00110001110" => rgb <= "010101";
when "00110001111" => rgb <= "011001";
when "00110010000" => rgb <= "010101";
when "00110010001" => rgb <= "011001";
when "00110010010" => rgb <= "010101";
when "00110010011" => rgb <= "010101";
when "00110100111" => rgb <= "010101";
when "00110101000" => rgb <= "010101";
when "00110101001" => rgb <= "011001";
when "00110101010" => rgb <= "011001";
when "00110101011" => rgb <= "011001";
when "00110101100" => rgb <= "011001";
when "00110101101" => rgb <= "010101";
when "00110101110" => rgb <= "011001";
when "00110101111" => rgb <= "011001";
when "00110110000" => rgb <= "011001";
when "00110110001" => rgb <= "011001";
when "00110110010" => rgb <= "010101";
when "00110110011" => rgb <= "010101";
when "00110110100" => rgb <= "010101";
when "00111000110" => rgb <= "010101";
when "00111000111" => rgb <= "000100";
when "00111001000" => rgb <= "010101";
when "00111001001" => rgb <= "011001";
when "00111001010" => rgb <= "011001";
when "00111001011" => rgb <= "011001";
when "00111001100" => rgb <= "011001";
when "00111001101" => rgb <= "011001";
when "00111001110" => rgb <= "011001";
when "00111001111" => rgb <= "011001";
when "00111010000" => rgb <= "011001";
when "00111010001" => rgb <= "011001";
when "00111010010" => rgb <= "011001";
when "00111010011" => rgb <= "010101";
when "00111010100" => rgb <= "000100";
when "00111010101" => rgb <= "010101";
when "00111100110" => rgb <= "010100";
when "00111100111" => rgb <= "010100";
when "00111101000" => rgb <= "010101";
when "00111101001" => rgb <= "011001";
when "00111101010" => rgb <= "011001";
when "00111101011" => rgb <= "011001";
when "00111101100" => rgb <= "011001";
when "00111101101" => rgb <= "011001";
when "00111101110" => rgb <= "011001";
when "00111101111" => rgb <= "011001";
when "00111110000" => rgb <= "011001";
when "00111110001" => rgb <= "011001";
when "00111110010" => rgb <= "011001";
when "00111110011" => rgb <= "010100";
when "00111110100" => rgb <= "000100";
when "00111110101" => rgb <= "010100";
when "01000000101" => rgb <= "010101";
when "01000000110" => rgb <= "010101";
when "01000000111" => rgb <= "010100";
when "01000001000" => rgb <= "010101";
when "01000001001" => rgb <= "011001";
when "01000001010" => rgb <= "011001";
when "01000001011" => rgb <= "011001";
when "01000001100" => rgb <= "011001";
when "01000001101" => rgb <= "010101";
when "01000001110" => rgb <= "011001";
when "01000001111" => rgb <= "011001";
when "01000010000" => rgb <= "011001";
when "01000010001" => rgb <= "011001";
when "01000010010" => rgb <= "010101";
when "01000010011" => rgb <= "010101";
when "01000010100" => rgb <= "010100";
when "01000010101" => rgb <= "010100";
when "01000010110" => rgb <= "010101";
when "01000100101" => rgb <= "010101";
when "01000100110" => rgb <= "010101";
when "01000100111" => rgb <= "000000";
when "01000101000" => rgb <= "010101";
when "01000101001" => rgb <= "010101";
when "01000101010" => rgb <= "010101";
when "01000101011" => rgb <= "010101";
when "01000101100" => rgb <= "010101";
when "01000101101" => rgb <= "010101";
when "01000101110" => rgb <= "010100";
when "01000101111" => rgb <= "010101";
when "01000110000" => rgb <= "010101";
when "01000110001" => rgb <= "010101";
when "01000110010" => rgb <= "010101";
when "01000110011" => rgb <= "010101";
when "01000110100" => rgb <= "000100";
when "01000110101" => rgb <= "010101";
when "01000110110" => rgb <= "010101";
when "01001000100" => rgb <= "010101";
when "01001000101" => rgb <= "000100";
when "01001000110" => rgb <= "000000";
when "01001000111" => rgb <= "000000";
when "01001001000" => rgb <= "010101";
when "01001001001" => rgb <= "010100";
when "01001001010" => rgb <= "010100";
when "01001001011" => rgb <= "010100";
when "01001001100" => rgb <= "011001";
when "01001001101" => rgb <= "011001";
when "01001001110" => rgb <= "011001";
when "01001001111" => rgb <= "011001";
when "01001010000" => rgb <= "010100";
when "01001010001" => rgb <= "010100";
when "01001010010" => rgb <= "010101";
when "01001010011" => rgb <= "010101";
when "01001010100" => rgb <= "000100";
when "01001010101" => rgb <= "010100";
when "01001010110" => rgb <= "010101";
when "01001100100" => rgb <= "010101";
when "01001100101" => rgb <= "010101";
when "01001100110" => rgb <= "000000";
when "01001101001" => rgb <= "010100";
when "01001101010" => rgb <= "010101";
when "01001101011" => rgb <= "011001";
when "01001101100" => rgb <= "011001";
when "01001101101" => rgb <= "011001";
when "01001101110" => rgb <= "010101";
when "01001101111" => rgb <= "011001";
when "01001110000" => rgb <= "011001";
when "01001110001" => rgb <= "010101";
when "01001110010" => rgb <= "010101";
when "01001110100" => rgb <= "010101";
when "01001110101" => rgb <= "000100";
when "01001110110" => rgb <= "010101";
when "01001110111" => rgb <= "100101";
when "01010000100" => rgb <= "010101";
when "01010000101" => rgb <= "010101";
when "01010000110" => rgb <= "010101";
when "01010001001" => rgb <= "010101";
when "01010001010" => rgb <= "010101";
when "01010001011" => rgb <= "010101";
when "01010001100" => rgb <= "011001";
when "01010001101" => rgb <= "011001";
when "01010001110" => rgb <= "011001";
when "01010001111" => rgb <= "011001";
when "01010010000" => rgb <= "010101";
when "01010010001" => rgb <= "010101";
when "01010010010" => rgb <= "010101";
when "01010010101" => rgb <= "000100";
when "01010010110" => rgb <= "010101";
when "01010010111" => rgb <= "010101";
when "01010100100" => rgb <= "010101";
when "01010100101" => rgb <= "010101";
when "01010100110" => rgb <= "010101";
when "01010101001" => rgb <= "011001";
when "01010101010" => rgb <= "010101";
when "01010101011" => rgb <= "010101";
when "01010101100" => rgb <= "011001";
when "01010101101" => rgb <= "011001";
when "01010101110" => rgb <= "011001";
when "01010101111" => rgb <= "011001";
when "01010110000" => rgb <= "010101";
when "01010110001" => rgb <= "011001";
when "01010110010" => rgb <= "010101";
when "01010110101" => rgb <= "010100";
when "01010110110" => rgb <= "010101";
when "01011000101" => rgb <= "010101";
when "01011000110" => rgb <= "000100";
when "01011001001" => rgb <= "010101";
when "01011001010" => rgb <= "010101";
when "01011001011" => rgb <= "010101";
when "01011001100" => rgb <= "011001";
when "01011001101" => rgb <= "011001";
when "01011001110" => rgb <= "011001";
when "01011001111" => rgb <= "011001";
when "01011010000" => rgb <= "010101";
when "01011010001" => rgb <= "011001";
when "01011010101" => rgb <= "010100";
when "01011010110" => rgb <= "010101";
when "01011100101" => rgb <= "010101";
when "01011100110" => rgb <= "000100";
when "01011101001" => rgb <= "010101";
when "01011101010" => rgb <= "011001";
when "01011101011" => rgb <= "011001";
when "01011101100" => rgb <= "011001";
when "01011101101" => rgb <= "011001";
when "01011101110" => rgb <= "011001";
when "01011101111" => rgb <= "010101";
when "01011110000" => rgb <= "010101";
when "01011110001" => rgb <= "010101";
when "01011110101" => rgb <= "010101";
when "01011110110" => rgb <= "010101";
when "01100000110" => rgb <= "010101";
when "01100001001" => rgb <= "010101";
when "01100001010" => rgb <= "010101";
when "01100001011" => rgb <= "010101";
when "01100001100" => rgb <= "011001";
when "01100001101" => rgb <= "011001";
when "01100001110" => rgb <= "011001";
when "01100001111" => rgb <= "011001";
when "01100010000" => rgb <= "011001";
when "01100010001" => rgb <= "010101";
when "01100010011" => rgb <= "101010";
when "01100010100" => rgb <= "101010";
when "01100010101" => rgb <= "011001";
when "01100100101" => rgb <= "101010";
when "01100100110" => rgb <= "101010";
when "01100100111" => rgb <= "101010";
when "01100101001" => rgb <= "000000";
when "01100101010" => rgb <= "000000";
when "01100101011" => rgb <= "010101";
when "01100101100" => rgb <= "010101";
when "01100101101" => rgb <= "010101";
when "01100101110" => rgb <= "010101";
when "01100101111" => rgb <= "010101";
when "01100110000" => rgb <= "000100";
when "01100110001" => rgb <= "000000";
when "01100110010" => rgb <= "010101";
when "01100110011" => rgb <= "101110";
when "01100110100" => rgb <= "101101";
when "01100110101" => rgb <= "101001";
when "01101000110" => rgb <= "101010";
when "01101000111" => rgb <= "101010";
when "01101001000" => rgb <= "010101";
when "01101001001" => rgb <= "000000";
when "01101001010" => rgb <= "000000";
when "01101001011" => rgb <= "000000";
when "01101001100" => rgb <= "000000";
when "01101001101" => rgb <= "000000";
when "01101001110" => rgb <= "000000";
when "01101001111" => rgb <= "000000";
when "01101010000" => rgb <= "000000";
when "01101010001" => rgb <= "000000";
when "01101010010" => rgb <= "010100";
when "01101010011" => rgb <= "101101";
when "01101010100" => rgb <= "101101";
when "01101010101" => rgb <= "101010";
when "01101100110" => rgb <= "101010";
when "01101100111" => rgb <= "010101";
when "01101101000" => rgb <= "000000";
when "01101101001" => rgb <= "000000";
when "01101101010" => rgb <= "000000";
when "01101101011" => rgb <= "000000";
when "01101101100" => rgb <= "000000";
when "01101101101" => rgb <= "000000";
when "01101101110" => rgb <= "000000";
when "01101101111" => rgb <= "000000";
when "01101110000" => rgb <= "000000";
when "01101110001" => rgb <= "000000";
when "01101110010" => rgb <= "000000";
when "01101110011" => rgb <= "011001";
when "01101110100" => rgb <= "101010";
when "01110000111" => rgb <= "010101";
when "01110001000" => rgb <= "000100";
when "01110001001" => rgb <= "000100";
when "01110001010" => rgb <= "000000";
when "01110001011" => rgb <= "000000";
when "01110001100" => rgb <= "000000";
when "01110001101" => rgb <= "000000";
when "01110001110" => rgb <= "000000";
when "01110001111" => rgb <= "000000";
when "01110010000" => rgb <= "000000";
when "01110010001" => rgb <= "000000";
when "01110010010" => rgb <= "000000";
when "01110010011" => rgb <= "010101";
when "01110100111" => rgb <= "010101";
when "01110101000" => rgb <= "011001";
when "01110101001" => rgb <= "011001";
when "01110101010" => rgb <= "010101";
when "01110101011" => rgb <= "010101";
when "01110101100" => rgb <= "010100";
when "01110101101" => rgb <= "000000";
when "01110101110" => rgb <= "000000";
when "01110101111" => rgb <= "000000";
when "01110110000" => rgb <= "000000";
when "01110110001" => rgb <= "000000";
when "01110110010" => rgb <= "010101";
when "01110110011" => rgb <= "010101";
when "01111000111" => rgb <= "010101";
when "01111001000" => rgb <= "010101";
when "01111001001" => rgb <= "011001";
when "01111001010" => rgb <= "011001";
when "01111001011" => rgb <= "010101";
when "01111001100" => rgb <= "010100";
when "01111001101" => rgb <= "100101";
when "01111001110" => rgb <= "010101";
when "01111001111" => rgb <= "010101";
when "01111010000" => rgb <= "010101";
when "01111010001" => rgb <= "011001";
when "01111010010" => rgb <= "010101";
when "01111010011" => rgb <= "010100";
when "01111010100" => rgb <= "010101";
when "01111101000" => rgb <= "010101";
when "01111101001" => rgb <= "010101";
when "01111101010" => rgb <= "011001";
when "01111101011" => rgb <= "010101";
when "01111101100" => rgb <= "010101";
when "01111101111" => rgb <= "010101";
when "01111110000" => rgb <= "010101";
when "01111110001" => rgb <= "011001";
when "01111110010" => rgb <= "011001";
when "01111110011" => rgb <= "010101";
when "10000001000" => rgb <= "010101";
when "10000001001" => rgb <= "010101";
when "10000001010" => rgb <= "011001";
when "10000001011" => rgb <= "010101";
when "10000001111" => rgb <= "100101";
when "10000010000" => rgb <= "010101";
when "10000010001" => rgb <= "010101";
when "10000010010" => rgb <= "010101";
when "10000010011" => rgb <= "010101";
when "10000101000" => rgb <= "010101";
when "10000101001" => rgb <= "010101";
when "10000101010" => rgb <= "010100";
when "10000101011" => rgb <= "010101";
when "10000110000" => rgb <= "010101";
when "10000110001" => rgb <= "010101";
when "10000110010" => rgb <= "010101";
when "10000110011" => rgb <= "010101";
when "10001001001" => rgb <= "010100";
when "10001001010" => rgb <= "010100";
when "10001001011" => rgb <= "010101";
when "10001010001" => rgb <= "010100";
when "10001010010" => rgb <= "010100";
when "10001010011" => rgb <= "010100";
when "10001010100" => rgb <= "010110";
when "10001101001" => rgb <= "010100";
when "10001101010" => rgb <= "010100";
when "10001101011" => rgb <= "010100";
when "10001110001" => rgb <= "010100";
when "10001110010" => rgb <= "010100";
when "10001110011" => rgb <= "010101";
when "10001110100" => rgb <= "010101";
when "10010001001" => rgb <= "010101";
when "10010001010" => rgb <= "010100";
when "10010001011" => rgb <= "010100";
when "10010001100" => rgb <= "010101";
when "10010010001" => rgb <= "010101";
when "10010010010" => rgb <= "010100";
when "10010010011" => rgb <= "010101";
when "10010010100" => rgb <= "010101";
when "10010101001" => rgb <= "010101";
when "10010101010" => rgb <= "010100";
when "10010101011" => rgb <= "010100";
when "10010101100" => rgb <= "010100";
when "10010110001" => rgb <= "010100";
when "10010110010" => rgb <= "010101";
when "10010110011" => rgb <= "010101";
when "10010110100" => rgb <= "010101";
when "10011001010" => rgb <= "010101";
when "10011001011" => rgb <= "010100";
when "10011001100" => rgb <= "010100";
when "10011010001" => rgb <= "010100";
when "10011010010" => rgb <= "010100";
when "10011010011" => rgb <= "010101";
when "10011101011" => rgb <= "010101";
when "10011101100" => rgb <= "010100";
when "10011110001" => rgb <= "010100";
when "10011110010" => rgb <= "010100";
when "10100001100" => rgb <= "010101";
when "10100010001" => rgb <= "010101";
when "10100010010" => rgb <= "010101";
when "10100101100" => rgb <= "010101";
when "10100101101" => rgb <= "011001";
when "10100110001" => rgb <= "010101";
when "10101001100" => rgb <= "011001";
when "10101001101" => rgb <= "011001";
when "10101010001" => rgb <= "011001";
when "10101101100" => rgb <= "011001";
when "10101101101" => rgb <= "011001";
when "10101110000" => rgb <= "010101";
when "10101110001" => rgb <= "011001";
when "10110001011" => rgb <= "101010";
when "10110001100" => rgb <= "011001";
when "10110001101" => rgb <= "011001";
when "10110010000" => rgb <= "010101";
when "10110010001" => rgb <= "011001";
when "10110010010" => rgb <= "101010";
when "10110101011" => rgb <= "101010";
when "10110101100" => rgb <= "011001";
when "10110101101" => rgb <= "011010";
when "10110110000" => rgb <= "011001";
when "10110110001" => rgb <= "011001";
when "10110110010" => rgb <= "101010";
when "10111010000" => rgb <= "010101";
when "10111010001" => rgb <= "011001";
when "10111010010" => rgb <= "101010";
when others => rgb <= "110011";



end case;

end if;

   end process;

   xy_address <= std_logic_vector(y_address) & std_logic_vector(x_address);
   
end;